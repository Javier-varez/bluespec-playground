package Zybo;

(* always_ready *)
interface Ifc_Top;
    (* prefix = "" *)
    method Bit#(4) led;
endinterface

endpackage
